module shift_add32
#(
	parameter WIDTH = 20
)
(
	input wire clk,rst,
	input wire signed[WIDTH-1:0] b0,
	input wire signed[WIDTH-1:0] b1,
	input wire signed[WIDTH-1:0] b2,
	input wire signed[WIDTH-1:0] b3,
	input wire signed[WIDTH-1:0] b4,
	input wire signed[WIDTH-1:0] b5,
	input wire signed[WIDTH-1:0] b6,
	input wire signed[WIDTH-1:0] b7,
	input wire signed[WIDTH-1:0] b8,
	input wire signed[WIDTH-1:0] b9,
	input wire signed[WIDTH-1:0] b10,
	input wire signed[WIDTH-1:0] b11,
	input wire signed[WIDTH-1:0] b12,
	input wire signed[WIDTH-1:0] b13,
	input wire signed[WIDTH-1:0] b14,
	input wire signed[WIDTH-1:0] b15,
	
	output reg signed[WIDTH-1:0] y1,
	output reg signed[WIDTH-1:0] y3,
	output reg signed[WIDTH-1:0] y5,
	output reg signed[WIDTH-1:0] y7,
	output reg signed[WIDTH-1:0] y9,
	output reg signed[WIDTH-1:0] y11,
	output reg signed[WIDTH-1:0] y13,
	output reg signed[WIDTH-1:0] y15,
	output reg signed[WIDTH-1:0] y17,
	output reg signed[WIDTH-1:0] y19,
	output reg signed[WIDTH-1:0] y21,
	output reg signed[WIDTH-1:0] y23,
	output reg signed[WIDTH-1:0] y25,
	output reg signed[WIDTH-1:0] y27,
	output reg signed[WIDTH-1:0] y29,
	output reg signed[WIDTH-1:0] y31
);

	wire signed [WIDTH-1:0] y1_d;
	wire signed [WIDTH-1:0] y3_d;
	wire signed [WIDTH-1:0] y5_d;
	wire signed [WIDTH-1:0] y7_d;
	wire signed [WIDTH-1:0] y9_d;
	wire signed [WIDTH-1:0] y11_d;
	wire signed [WIDTH-1:0] y13_d;
	wire signed [WIDTH-1:0] y15_d;
	wire signed [WIDTH-1:0] y17_d;
	wire signed [WIDTH-1:0] y19_d;
	wire signed [WIDTH-1:0] y21_d;
	wire signed [WIDTH-1:0] y23_d;
	wire signed [WIDTH-1:0] y25_d;
	wire signed [WIDTH-1:0] y27_d;
	wire signed [WIDTH-1:0] y29_d;
	wire signed [WIDTH-1:0] y31_d;
	
	always @ (posedge clk)
	begin
//		if(!rst_b) begin
		if(rst) begin
				y1 <= 0;
				y3 <= 0;
				y5 <= 0;
				y7 <= 0;
				y9 <= 0;
				y11 <= 0;
				y13 <= 0;
				y15 <= 0;
				y17 <= 0;
				y19 <= 0;
				y21 <= 0;
				y23 <= 0;
				y25 <= 0;
				y27 <= 0;
				y29 <= 0;
				y31 <= 0;
		end
		else begin
				y1 <= y1_d;
				y3 <= y3_d;
				y5 <= y5_d;
				y7 <= y7_d;
				y9 <= y9_d;
				y11 <= y11_d;
				y13 <= y13_d;
				y15 <= y15_d;
				y17 <= y17_d;
				y19 <= y19_d;
				y21 <= y21_d;
				y23 <= y23_d;
				y25 <= y25_d;
				y27 <= y27_d;
				y29 <= y29_d;
				y31 <= y31_d;
				
		end
	end
	
	assign y1_d = {b0,1'b0}+{b0,3'b000}+{b0,4'b0000}+{b0,6'b000000}+{b1,1'b0}+{b1,3'b000}+{b1,4'b0000}+{b1,6'b000000}+{b2,3'b000}+{b2,4'b0000}+{b2,6'b000000}+b3+{b3,2'b00}+{b3,4'b0000}+{b3,6'b000000}+{b4,1'b0}+{b4,4'b0000}+{b4,6'b000000}+{b5,1'b0}+{b5,2'b00}+{b5,3'b000}+{b5,6'b000000}+b6+{b6,3'b000}+{b6,6'b000000}+b7+{b7,1'b0}+{b7,6'b000000}+b8+{b8,2'b00}+{b8,3'b000}+{b8,4'b0000}+{b8,5'b00000}+{b9,1'b0}+{b9,2'b00}+{b9,4'b0000}+{b9,5'b00000}+{b10,1'b0}+{b10,2'b00}+{b10,3'b000}+{b10,5'b00000}+{b11,1'b0}+{b11,2'b00}+{b11,5'b00000}+b12+{b12,1'b0}+{b12,2'b00}+{b12,3'b000}+{b12,4'b0000}+{b13,1'b0}+{b13,2'b00}+{b13,4'b0000}+b14+{b14,2'b00}+{b14,3'b000}+{b15,2'b00};

	assign y3_d = {b0,1'b0}+{b0,3'b000}+{b0,4'b0000}+{b0,6'b000000}+{b1,1'b0}+{b1,4'b0000}+{b1,6'b000000}+b2+{b2,1'b0}+{b2,6'b000000}+{b3,1'b0}+{b3,2'b00}+{b3,3'b000}+{b3,5'b00000}+{b4,1'b0}+{b4,2'b00}+{b4,4'b0000}-{b5,2'b00}-b6-{b6,1'b0}-{b6,2'b00}-{b6,3'b000}-{b6,4'b0000}-{b7,1'b0}-{b7,2'b00}-{b7,4'b0000}-{b7,5'b00000}-b8-{b8,3'b000}-{b8,6'b000000}-b9-{b9,2'b00}-{b9,4'b0000}-{b9,6'b000000}-{b10,1'b0}-{b10,3'b000}-{b10,4'b0000}-{b10,6'b000000}-{b11,3'b000}-{b11,4'b0000}-{b11,6'b000000}-{b12,1'b0}-{b12,2'b00}-{b12,3'b000}-{b12,6'b000000}-b13-{b13,2'b00}-{b13,3'b000}-{b13,4'b0000}-{b13,5'b00000}-{b14,1'b0}-{b14,2'b00}-{b14,5'b00000}-b15-{b15,2'b00}-{b15,3'b000};

	assign y5_d = {b0,3'b000}+{b0,4'b0000}+{b0,6'b000000}+b1+{b1,1'b0}+{b1,6'b000000}+b2+{b2,1'b0}+{b2,2'b00}+{b2,3'b000}+{b2,4'b0000}-b3-{b3,2'b00}-{b3,3'b000}-{b4,1'b0}-{b4,2'b00}-{b4,4'b0000}-{b4,5'b00000}-{b5,1'b0}-{b5,4'b0000}-{b5,6'b000000}-{b6,1'b0}-{b6,3'b000}-{b6,4'b0000}-{b6,6'b000000}-{b7,1'b0}-{b7,2'b00}-{b7,3'b000}-{b7,6'b000000}-{b8,1'b0}-{b8,2'b00}-{b8,3'b000}-{b8,5'b00000}-{b9,2'b00}+{b10,1'b0}+{b10,2'b00}+{b10,5'b00000}+b11+{b11,3'b000}+{b11,6'b000000}+{b12,1'b0}+{b12,3'b000}+{b12,4'b0000}+{b12,6'b000000}+b13+{b13,2'b00}+{b13,4'b0000}+{b13,6'b000000}+b14+{b14,2'b00}+{b14,3'b000}+{b14,4'b0000}+{b14,5'b00000}+{b15,1'b0}+{b15,2'b00}+{b15,4'b0000};

	assign y7_d = b0+{b0,2'b00}+{b0,4'b0000}+{b0,6'b000000}+{b1,1'b0}+{b1,2'b00}+{b1,3'b000}+{b1,5'b00000}-b2-{b2,2'b00}-{b2,3'b000}-b3-{b3,1'b0}-{b3,6'b000000}-{b4,1'b0}-{b4,3'b000}-{b4,4'b0000}-{b4,6'b000000}-b5-{b5,3'b000}-{b5,6'b000000}-{b6,1'b0}-{b6,2'b00}-{b6,4'b0000}+{b7,1'b0}+{b7,2'b00}+{b7,5'b00000}+{b8,1'b0}+{b8,4'b0000}+{b8,6'b000000}+{b9,3'b000}+{b9,4'b0000}+{b9,6'b000000}+{b10,1'b0}+{b10,2'b00}+{b10,4'b0000}+{b10,5'b00000}-{b11,2'b00}-b12-{b12,2'b00}-{b12,3'b000}-{b12,4'b0000}-{b12,5'b00000}-{b13,1'b0}-{b13,3'b000}-{b13,4'b0000}-{b13,6'b000000}-{b14,1'b0}-{b14,2'b00}-{b14,3'b000}-{b14,6'b000000}-b15-{b15,1'b0}-{b15,2'b00}-{b15,3'b000}-{b15,4'b0000};

	assign y9_d = {b0,1'b0}+{b0,4'b0000}+{b0,6'b000000}+{b1,1'b0}+{b1,2'b00}+{b1,4'b0000}-{b2,1'b0}-{b2,2'b00}-{b2,4'b0000}-{b2,5'b00000}-{b3,1'b0}-{b3,3'b000}-{b3,4'b0000}-{b3,6'b000000}-b4-{b4,2'b00}-{b4,3'b000}-{b4,4'b0000}-{b4,5'b00000}+b5+{b5,1'b0}+{b5,2'b00}+{b5,3'b000}+{b5,4'b0000}+{b6,1'b0}+{b6,2'b00}+{b6,3'b000}+{b6,6'b000000}+b7+{b7,2'b00}+{b7,4'b0000}+{b7,6'b000000}+b8+{b8,1'b0}+{b8,2'b00}+{b8,3'b000}+{b8,4'b0000}-{b9,1'b0}-{b9,2'b00}-{b9,3'b000}-{b9,5'b00000}-{b10,1'b0}-{b10,3'b000}-{b10,4'b0000}-{b10,6'b000000}-b11-{b11,1'b0}-{b11,6'b000000}+{b12,2'b00}+b13+{b13,3'b000}+{b13,6'b000000}+{b14,3'b000}+{b14,4'b0000}+{b14,6'b000000}+{b15,1'b0}+{b15,2'b00}+{b15,5'b00000};

	assign y11_d = {b0,1'b0}+{b0,2'b00}+{b0,3'b000}+{b0,6'b000000}-{b1,2'b00}-{b2,1'b0}-{b2,4'b0000}-{b2,6'b000000}-b3-{b3,3'b000}-{b3,6'b000000}+b4+{b4,2'b00}+{b4,3'b000}+b5+{b5,2'b00}+{b5,4'b0000}+{b5,6'b000000}+b6+{b6,1'b0}+{b6,6'b000000}-{b7,1'b0}-{b7,2'b00}-{b7,4'b0000}-{b8,3'b000}-{b8,4'b0000}-{b8,6'b000000}-b9-{b9,2'b00}-{b9,3'b000}-{b9,4'b0000}-{b9,5'b00000}+b10+{b10,1'b0}+{b10,2'b00}+{b10,3'b000}+{b10,4'b0000}+{b11,1'b0}+{b11,3'b000}+{b11,4'b0000}+{b11,6'b000000}+{b12,1'b0}+{b12,2'b00}+{b12,4'b0000}+{b12,5'b00000}-{b13,1'b0}-{b13,2'b00}-{b13,5'b00000}-{b14,1'b0}-{b14,3'b000}-{b14,4'b0000}-{b14,6'b000000}-{b15,1'b0}-{b15,2'b00}-{b15,3'b000}-{b15,5'b00000};

	assign y13_d = b0+{b0,3'b000}+{b0,6'b000000}-b1-{b1,1'b0}-{b1,2'b00}-{b1,3'b000}-{b1,4'b0000}-{b2,1'b0}-{b2,3'b000}-{b2,4'b0000}-{b2,6'b000000}-{b3,1'b0}-{b3,2'b00}-{b3,4'b0000}+{b4,1'b0}+{b4,2'b00}+{b4,3'b000}+{b4,6'b000000}+b5+{b5,1'b0}+{b5,6'b000000}-{b6,1'b0}-{b6,2'b00}-{b6,5'b00000}-{b7,1'b0}-{b7,3'b000}-{b7,4'b0000}-{b7,6'b000000}-b8-{b8,2'b00}-{b8,3'b000}+{b9,1'b0}+{b9,4'b0000}+{b9,6'b000000}+b10+{b10,2'b00}+{b10,3'b000}+{b10,4'b0000}+{b10,5'b00000}-{b11,1'b0}-{b11,2'b00}-{b11,3'b000}-{b11,5'b00000}-{b12,3'b000}-{b12,4'b0000}-{b12,6'b000000}-{b13,2'b00}+b14+{b14,2'b00}+{b14,4'b0000}+{b14,6'b000000}+{b15,1'b0}+{b15,2'b00}+{b15,4'b0000}+{b15,5'b00000};

	assign y15_d = b0+{b0,1'b0}+{b0,6'b000000}-{b1,1'b0}-{b1,2'b00}-{b1,4'b0000}-{b1,5'b00000}-{b2,1'b0}-{b2,2'b00}-{b2,3'b000}-{b2,6'b000000}+{b3,1'b0}+{b3,2'b00}+{b3,5'b00000}+b4+{b4,2'b00}+{b4,4'b0000}+{b4,6'b000000}-{b5,1'b0}-{b5,2'b00}-{b5,4'b0000}-{b6,1'b0}-{b6,3'b000}-{b6,4'b0000}-{b6,6'b000000}+{b7,2'b00}+{b8,1'b0}+{b8,3'b000}+{b8,4'b0000}+{b8,6'b000000}+b9+{b9,2'b00}+{b9,3'b000}-{b10,3'b000}-{b10,4'b0000}-{b10,6'b000000}-b11-{b11,1'b0}-{b11,2'b00}-{b11,3'b000}-{b11,4'b0000}+{b12,1'b0}+{b12,4'b0000}+{b12,6'b000000}+{b13,1'b0}+{b13,2'b00}+{b13,3'b000}+{b13,5'b00000}-b14-{b14,3'b000}-{b14,6'b000000}-b15-{b15,2'b00}-{b15,3'b000}-{b15,4'b0000}-{b15,5'b00000};

	assign y17_d = b0+{b0,2'b00}+{b0,3'b000}+{b0,4'b0000}+{b0,5'b00000}-b1-{b1,3'b000}-{b1,6'b000000}-{b2,1'b0}-{b2,2'b00}-{b2,3'b000}-{b2,5'b00000}+{b3,1'b0}+{b3,4'b0000}+{b3,6'b000000}+b4+{b4,1'b0}+{b4,2'b00}+{b4,3'b000}+{b4,4'b0000}-{b5,3'b000}-{b5,4'b0000}-{b5,6'b000000}-b6-{b6,2'b00}-{b6,3'b000}+{b7,1'b0}+{b7,3'b000}+{b7,4'b0000}+{b7,6'b000000}-{b8,2'b00}-{b9,1'b0}-{b9,3'b000}-{b9,4'b0000}-{b9,6'b000000}+{b10,1'b0}+{b10,2'b00}+{b10,4'b0000}+b11+{b11,2'b00}+{b11,4'b0000}+{b11,6'b000000}-{b12,1'b0}-{b12,2'b00}-{b12,5'b00000}-{b13,1'b0}-{b13,2'b00}-{b13,3'b000}-{b13,6'b000000}+{b14,1'b0}+{b14,2'b00}+{b14,4'b0000}+{b14,5'b00000}+b15+{b15,1'b0}+{b15,6'b000000};

	assign y19_d = {b0,1'b0}+{b0,2'b00}+{b0,4'b0000}+{b0,5'b00000}-b1-{b1,2'b00}-{b1,4'b0000}-{b1,6'b000000}-{b2,2'b00}+{b3,3'b000}+{b3,4'b0000}+{b3,6'b000000}-{b4,1'b0}-{b4,2'b00}-{b4,3'b000}-{b4,5'b00000}-b5-{b5,2'b00}-{b5,3'b000}-{b5,4'b0000}-{b5,5'b00000}+{b6,1'b0}+{b6,4'b0000}+{b6,6'b000000}+b7+{b7,2'b00}+{b7,3'b000}-{b8,1'b0}-{b8,3'b000}-{b8,4'b0000}-{b8,6'b000000}+{b9,1'b0}+{b9,2'b00}+{b9,5'b00000}+b10+{b10,1'b0}+{b10,6'b000000}-{b11,1'b0}-{b11,2'b00}-{b11,3'b000}-{b11,6'b000000}-{b12,1'b0}-{b12,2'b00}-{b12,4'b0000}+{b13,1'b0}+{b13,3'b000}+{b13,4'b0000}+{b13,6'b000000}-b14-{b14,1'b0}-{b14,2'b00}-{b14,3'b000}-{b14,4'b0000}-b15-{b15,3'b000}-{b15,6'b000000};

	assign y21_d = {b0,1'b0}+{b0,2'b00}+{b0,3'b000}+{b0,5'b00000}-{b1,1'b0}-{b1,3'b000}-{b1,4'b0000}-{b1,6'b000000}+{b2,1'b0}+{b2,2'b00}+{b2,5'b00000}+{b3,1'b0}+{b3,2'b00}+{b3,4'b0000}+{b3,5'b00000}-{b4,1'b0}-{b4,3'b000}-{b4,4'b0000}-{b4,6'b000000}+b5+{b5,1'b0}+{b5,2'b00}+{b5,3'b000}+{b5,4'b0000}+b6+{b6,2'b00}+{b6,3'b000}+{b6,4'b0000}+{b6,5'b00000}-{b7,3'b000}-{b7,4'b0000}-{b7,6'b000000}+{b8,1'b0}+{b8,2'b00}+{b8,4'b0000}+b9+{b9,1'b0}+{b9,6'b000000}-b10-{b10,2'b00}-{b10,4'b0000}-{b10,6'b000000}+b11+{b11,2'b00}+{b11,3'b000}+b12+{b12,3'b000}+{b12,6'b000000}-{b13,1'b0}-{b13,4'b0000}-{b13,6'b000000}+{b14,2'b00}+{b15,1'b0}+{b15,2'b00}+{b15,3'b000}+{b15,6'b000000};

	assign y23_d = {b0,1'b0}+{b0,2'b00}+{b0,5'b00000}-{b1,3'b000}-{b1,4'b0000}-{b1,6'b000000}+b2+{b2,3'b000}+{b2,6'b000000}-{b3,2'b00}-b4-{b4,1'b0}-{b4,6'b000000}+{b5,1'b0}+{b5,3'b000}+{b5,4'b0000}+{b5,6'b000000}-{b6,1'b0}-{b6,2'b00}-{b6,3'b000}-{b6,5'b00000}-b7-{b7,1'b0}-{b7,2'b00}-{b7,3'b000}-{b7,4'b0000}+b8+{b8,2'b00}+{b8,4'b0000}+{b8,6'b000000}-{b9,1'b0}-{b9,2'b00}-{b9,3'b000}-{b9,6'b000000}+b10+{b10,2'b00}+{b10,3'b000}+b11+{b11,2'b00}+{b11,3'b000}+{b11,4'b0000}+{b11,5'b00000}-{b12,1'b0}-{b12,3'b000}-{b12,4'b0000}-{b12,6'b000000}+{b13,1'b0}+{b13,2'b00}+{b13,4'b0000}+{b13,5'b00000}+{b14,1'b0}+{b14,2'b00}+{b14,4'b0000}-{b15,1'b0}-{b15,4'b0000}-{b15,6'b000000};

	assign y25_d = b0+{b0,1'b0}+{b0,2'b00}+{b0,3'b000}+{b0,4'b0000}-{b1,1'b0}-{b1,2'b00}-{b1,3'b000}-{b1,6'b000000}+{b2,1'b0}+{b2,3'b000}+{b2,4'b0000}+{b2,6'b000000}-b3-{b3,2'b00}-{b3,3'b000}-{b3,4'b0000}-{b3,5'b00000}+{b4,2'b00}+{b5,1'b0}+{b5,2'b00}+{b5,4'b0000}+{b5,5'b00000}-{b6,3'b000}-{b6,4'b0000}-{b6,6'b000000}+{b7,1'b0}+{b7,4'b0000}+{b7,6'b000000}-{b8,1'b0}-{b8,2'b00}-{b8,5'b00000}-{b9,1'b0}-{b9,2'b00}-{b9,4'b0000}+b10+{b10,3'b000}+{b10,6'b000000}-{b11,1'b0}-{b11,3'b000}-{b11,4'b0000}-{b11,6'b000000}+b12+{b12,1'b0}+{b12,6'b000000}-b13-{b13,2'b00}-{b13,3'b000}-{b14,1'b0}-{b14,2'b00}-{b14,3'b000}-{b14,5'b00000}+b15+{b15,2'b00}+{b15,4'b0000}+{b15,6'b000000};

	assign y27_d = {b0,1'b0}+{b0,2'b00}+{b0,4'b0000}-b1-{b1,2'b00}-{b1,3'b000}-{b1,4'b0000}-{b1,5'b00000}+b2+{b2,2'b00}+{b2,4'b0000}+{b2,6'b000000}-{b3,1'b0}-{b3,3'b000}-{b3,4'b0000}-{b3,6'b000000}+b4+{b4,3'b000}+{b4,6'b000000}-{b5,1'b0}-{b5,2'b00}-{b5,5'b00000}-{b6,2'b00}+{b7,1'b0}+{b7,2'b00}+{b7,3'b000}+{b7,5'b00000}-{b8,1'b0}-{b8,2'b00}-{b8,3'b000}-{b8,6'b000000}+{b9,1'b0}+{b9,3'b000}+{b9,4'b0000}+{b9,6'b000000}-{b10,1'b0}-{b10,4'b0000}-{b10,6'b000000}+{b11,1'b0}+{b11,2'b00}+{b11,4'b0000}+{b11,5'b00000}-b12-{b12,2'b00}-{b12,3'b000}-b13-{b13,1'b0}-{b13,2'b00}-{b13,3'b000}-{b13,4'b0000}+b14+{b14,1'b0}+{b14,6'b000000}-{b15,3'b000}-{b15,4'b0000}-{b15,6'b000000};

	assign y29_d = b0+{b0,2'b00}+{b0,3'b000}-{b1,1'b0}-{b1,2'b00}-{b1,5'b00000}+b2+{b2,2'b00}+{b2,3'b000}+{b2,4'b0000}+{b2,5'b00000}-{b3,1'b0}-{b3,2'b00}-{b3,3'b000}-{b3,6'b000000}+{b4,3'b000}+{b4,4'b0000}+{b4,6'b000000}-{b5,1'b0}-{b5,3'b000}-{b5,4'b0000}-{b5,6'b000000}+b6+{b6,2'b00}+{b6,4'b0000}+{b6,6'b000000}-b7-{b7,3'b000}-{b7,6'b000000}+{b8,1'b0}+{b8,2'b00}+{b8,4'b0000}+{b8,5'b00000}-b9-{b9,1'b0}-{b9,2'b00}-{b9,3'b000}-{b9,4'b0000}+{b10,2'b00}+{b11,1'b0}+{b11,2'b00}+{b11,4'b0000}-{b12,1'b0}-{b12,2'b00}-{b12,3'b000}-{b12,5'b00000}+b13+{b13,1'b0}+{b13,6'b000000}-{b14,1'b0}-{b14,4'b0000}-{b14,6'b000000}+{b15,1'b0}+{b15,3'b000}+{b15,4'b0000}+{b15,6'b000000};

	assign y31_d = {b0,2'b00}-b1-{b1,2'b00}-{b1,3'b000}+{b2,1'b0}+{b2,2'b00}+{b2,4'b0000}-b3-{b3,1'b0}-{b3,2'b00}-{b3,3'b000}-{b3,4'b0000}+{b4,1'b0}+{b4,2'b00}+{b4,5'b00000}-{b5,1'b0}-{b5,2'b00}-{b5,3'b000}-{b5,5'b00000}+{b6,1'b0}+{b6,2'b00}+{b6,4'b0000}+{b6,5'b00000}-b7-{b7,2'b00}-{b7,3'b000}-{b7,4'b0000}-{b7,5'b00000}+b8+{b8,1'b0}+{b8,6'b000000}-b9-{b9,3'b000}-{b9,6'b000000}+{b10,1'b0}+{b10,2'b00}+{b10,3'b000}+{b10,6'b000000}-{b11,1'b0}-{b11,4'b0000}-{b11,6'b000000}+b12+{b12,2'b00}+{b12,4'b0000}+{b12,6'b000000}-{b13,3'b000}-{b13,4'b0000}-{b13,6'b000000}+{b14,1'b0}+{b14,3'b000}+{b14,4'b0000}+{b14,6'b000000}-{b15,1'b0}-{b15,3'b000}-{b15,4'b0000}-{b15,6'b000000};
	
	//x90 = {b0,6'b000000} + {b0,4'b0000} + {b0,3'b000} + {b0,1'b0}
	//x88 = {b0,6'b000000} + {b0,4'b0000} + {b0,3'b000}
	//x87 = {b0,6'b000000} + {b0,4'b0000} + {b0,2'b00} + {b0,1'b0} + b0
	//x85 = {b0,6'b000000} + {b0,4'b0000} + {b0,2'b00} + b0
	//x82 = {b0,6'b000000} + {b0,4'b0000} + {b0,1'b0}
	//x80 = {b0,6'b000000} + {b0,4'b0000} 
	//x78 = {b0,6'b000000} + {b0,3'b000} + {b0,2'b00} + {b0,1'b0}
	//x73 = {b0,6'b000000} + {b0,3'b000} + b0
	//x70 = {b0,6'b000000} + {b0,2'b00} + {b0,1'b0}
	//x67 = {b0,6'b000000} + {b0,1'b0} + b0
	//x61 = {b0,5'b00000} + {b0,4'b0000} + {b0,3'b000} + {b0,2'b00} + b0
	//x57 = {b0,5'b00000} + {b0,4'b0000} + {b0,3'b000} + {b0,1'b0}
	//x54 = {b0,5'b00000} + {b0,4'b0000} + {b0,2'b00} + {b0,1'b0}
	//x46 = {b0,5'b00000} + {b0,3'b000} + {b0,2'b00} + {b0,1'b0}
	//x43 = {b0,5'b00000} + {b0,3'b000} + {b0,1'b0} + b0
	//x38 = {b0,5'b00000} + {b0,2'b00} + {b0,1'b0}
	//x31 = {b0,4'b0000} + {b0,3'b000} + {b0,2'b00} + {b0,1'b0} + b0
	//x25 = {b0,4'b0000} + {b0,3'b000} + {b0,1'b0}
	//x22 = {b0,4'b0000} + {b0,2'b00} + {b0,1'b0}
	//x13 = {b0,3'b000} + {b0,2'b00} + b0
	//x9  = {b0,3'b000} + {b0,1'b0}
	//x4  = {b0,2'b00}
	
	
endmodule 